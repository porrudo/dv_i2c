`include "base_test.sv"

`include "test_dummy.sv"
`include "test_reset.sv"
`include "test_write.sv"
//other tests